
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package CORDIC_package is 
    
    TYPE state IS
        (ST0,ST1,ST2,ST3,ST4,ST5,ST6,ST7);
            
end package CORDIC_package;